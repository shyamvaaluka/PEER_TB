//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//	version					:	0.1
//	file name				: ecc.sv
//	description			:	This module includes the encrypter and decrypter designs for both of the ports. Simply, it instantiates the encrypter design for
//										both the ports and connects the recieved inputs to it and produce the encrypted data as outputs. In a similar, this design will
//										recieve the encrypted (whether it might be corrected or error freee) and the decrypter designs will outputs the decrypted data
//										as output.
//										
//	parametrs used	:	DATA_WIDTH	=	8 ->	This parameter defines the data width of input data and accordingly the data width of the output will be
//																				calculated it self.
// 
//  Input Ports   	:	i_data_a,i_data_b		:	This is the input pin to the design and once the change happened in this port automatically the encrypted
//  																				data will	be caluclated by passing to the respective encrypted design.
//										i_enc_dina,					:	These are input pins (which is nothing but encrypted read data) and this will be connected to input pins
//										i_enc_dinb						of the data decrypter design's.
//										
//
//  Output Ports		:	o_enc_data_a,				: These are the output port of this module, this ports will be used to collect the encrypted outputs from the
//  									o_enc_data_b					data encrypter desing's.
//										o_decr_data_a,			:	These are the output port of this module, this ports will be used to collect the decrypted data generated by
//										o_decr_data_b					the data decrypter design's.
//										o_errora,o_errorb		:	These are the output ports of this module,this ports will be connected with the errror out ports of each
//																					data decrypter design's error output ports.
//
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module ecc #(parameter DATA_WIDTH = 8)
						(	input 	[DATA_WIDTH-1												:0]	i_data_a,
							input 	[DATA_WIDTH-1												:0]	i_data_b,
							input 	[DATA_WIDTH + $clog2(DATA_WIDTH) +1	:0]	i_enc_dina,
							input 	[DATA_WIDTH + $clog2(DATA_WIDTH) +1	:0]	i_enc_dinb,
							output 	[DATA_WIDTH + $clog2(DATA_WIDTH) +1	:0]	o_enc_data_a,
							output 	[DATA_WIDTH + $clog2(DATA_WIDTH) +1	:0]	o_enc_data_b,
							output 	[DATA_WIDTH - 1										 	:0]	o_decr_data_a,
							output 	[DATA_WIDTH - 1										 	:0]	o_decr_data_b,
							output	                                      	o_errora,
							output	                                      	o_errorb
						);
		
		//Encrypter and Decrypter Design's instantiation's
		hamming_encoder			#(DATA_WIDTH)	ENC_DUTA		(	.i_data(i_data_a),
									 																	.o_enc_data(o_enc_data_a));
		hamming_encoder			#(DATA_WIDTH)	ENC_DUTB		(	.i_data(i_data_b),
																										.o_enc_data(o_enc_data_b));
		hamming_decoder			#(DATA_WIDTH)	DE_ENC_DUTA	(	.i_enc_data(i_enc_dina),
							 		 																	.o_error(o_errora),
							 		 																	.o_decr_data(o_decr_data_a));
		hamming_decoder			#(DATA_WIDTH)	DE_ENC_DUTB	(	.i_enc_data(i_enc_dinb),
																										.o_error(o_errorb),
																										.o_decr_data(o_decr_data_b));

endmodule : ecc
